module ControllerHours
(
    input clk,
)

    reg[0:3] curr_state;
    reg[0:3] next_state;

    always @(*)
    begin
        case(curr_state)
    end
        